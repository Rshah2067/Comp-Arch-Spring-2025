//For R type instructions needs to distinguish which ALU module is being used